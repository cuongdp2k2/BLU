parameter Q = 8380417 ;  