module NTT #(
    parameter DATA_WIDTH = 8 ,
    parameter DATA_NUM   = 8 
) (
    input logic clk_i , reset_ni ,
    input logic [DATA_WIDTH-1:0] data_i [DATA_NUM-1:0],

    output
);
endmodule : NTT 